`timescale 10ns/1ns
module MIPS_test;
reg clk,reset;

initial 
begin
	clk=0;
end

endmodule
