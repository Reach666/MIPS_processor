module adder_30(C,A,B);

input A,B;
output C;

wire [29:0]A,B,C;

assign C = A + B;

endmodule 